module top();

dut u_dut();
router u_router();

endmodule
